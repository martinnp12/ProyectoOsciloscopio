----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 19.05.2021 09:34:11
-- Design Name: 
-- Module Name: CharacterROM - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.oscilloscope_pkg.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CharacterROM is
    Port ( clk_i : in STD_LOGIC;
           reset_i : in STD_LOGIC;
           addr_i : in STD_LOGIC_VECTOR (7 downto 0);
           data_o : out STD_LOGIC_VECTOR (7 downto 0));
end CharacterROM;

architecture Behavioral of CharacterROM is
  signal rom : character_rom_t := (
  -- 0: code x00
   "00111100",    
   "01100110",
   "01100110",
   "01100110",
   "01100110",
   "01100110",
   "01100110",
   "00111100",
   -- 1: code x01
   "00011100", 
   "00111100",
   "01101100",
   "00001100",
   "00001100",
   "00001100",
   "00001100",
   -- 2 : code x02
   "00111111",   
   "00111100",
   "01100110",
   "01100110",
   "00001100",
   "00011000",
   "00110000",
   "01100000",
   "01111110",   
   -- 3 : code x03
   "00111100", 
   "01100110",
   "00000110",
   "00011100",
   "00000110",
   "00000110",
   "01100110",
   "00111100", 
   -- 4 code x04
   "00011100",   
   "00111100",
   "01101100",
   "11001100",
   "11111111",
   "00001100",
   "00001100",
   "00001100",
   -- 5: code x05
   "01111110",    
   "01100000",
   "01100000",
   "01111100",
   "00000110",
   "00000011",
   "01100110",
   "00111100",
   -- 6 code x06
   "00111100",   
   "01100110",
   "01100110",
   "01100000",
   "01111100",
   "01100010",
   "00110110",
   "00011100",
   -- 7 code x07
   "01111110",   
   "01100110",
   "00001100",
   "00011000",
   "00110000",
   "00110000",
   "00110000",
   "00110000",   
   -- 8 code x08
   "00111100",
   "01100110",
   "01100110",
   "00111100",
   "00111100",
   "01100110",
   "01100110",
   "00111100", 
     -- 9 code x09
   "00111100",
   "01100110",
   "01100110",
   "00111110",
   "00000110",
   "01100110",
   "01100110",
   "00111100",
   -- . code x0A
   "00000000", 
   "00000000",
   "00000000",
   "00000000",
   "00000000",
   "00000000",
   "00110000",
   "00110000", 
   --: code x0B
   "00000000", 
   "00000000",
   "00000000",
   "00110000",
   "00110000",
   "00000000",
   "00110000",
   "00110000",
   -- = code x0C
   "00000000", 
   "01111110",
   "01111110",
   "00000000",
   "00000000",
   "01111110",
   "01111110",
   "00000000",
   -- u code x0D
   "00000000", 
   "00000000",
   "00000000",
   "00100010",
   "00100010",
   "00100010",
   "00100110",
   "00011010",
   -- m code x0E
   "00000000", 
   "00000000",
   "01101110",
   "10010001",
   "10010001",
   "10010001",
   "10010001",
   "10010001",
   -- V code x0F
   "10000001", 
   "10000001",
   "01000010",
   "01000010",
   "00100100",
   "00100100",
   "00011000",
   "00011000",
   -- s code x10
   "00000000", 
   "00000000",
   "00111000",
   "01000000",
   "00111000",
   "00000100",
   "01000100",
   "00111000",
   -- / code x11
   "00000010", 
   "00000110",
   "00001100",
   "00011000",
   "00110000",
   "01100000",
   "01000000",
   "10000000",
   -- A code x12
   "00011000", 
   "00100100",
   "01000010",
   "01000010",
   "01111110",
   "01000010",
   "01000010",
   "01000010",
   --U code x13
   "01000010", 
   "01000010",
   "01000010",
   "01000010",
   "01000010",
   "01000010",
   "00100100",
   "00011000",
   --T code x14
   "11111110", 
   "00010000",
   "00010000",
   "00010000",
   "00010000",
   "00010000",
   "00010000",
   "00010000",
   --O code x15
   "00111100", 
   "01000010",
   "10000001",
   "10000001",
   "10000001",
   "10000001",
   "01000010",
   "00111100",
   -- NULL code x16
   "00000000", 
   "00000000",
   "00000000",
   "00000000",
   "00000000",
   "00000000",
   "00000000",
   "00000000",
   -- x code x17
   "00000000", 
   "00000000",
   "01100011",
   "00110110",
   "00011100",
   "00011100",
   "00110110",
   "01100011",
   -- i code x18
   "00000000", 
   "00001100",
   "00001100",
   "00000000",
   "00001100",
   "00001100",
   "00001100",
   "00001100",
   -- n code x18
   "00000000", 
   "00000000",
   "00000000",
   "00000000",
   "00001110",
   "00010001",
   "00010001",
   "00010001",
   -- - code x19
   "00000000", 
   "00000000",
   "00000000",
   "01111110",
   "01111110",
   "00000000",
   "00000000",
   "00000000",
   -- p code x1A
   "00000000", 
   "00000000",
   "00010110",
   "00011001",
   "00010001",
   "00011110",
   "00010000",
   "00010000",
   -- a code x1B
   "00000000", 
   "00000000",
   "00000000",
   "00001110",
   "00000001",
   "00001111",
   "00010001",
   "00001111",
   -- v code x1C
   "00000000", 
   "00000000",
   "00000000",
   "00010001",
   "00010001",
   "00010001",
   "00001010",
   "00000100",
   -- g code x1D
   "00000000", 
   "00001111",
   "00001111",
   "00010001",
   "00010001",
   "00001111",
   "00000001",
   "00011110", 
   -- k code x1E
   "00000000",
   "00001000",
   "00001000",
   "00001001",
   "00001010",
   "00001100",
   "00001010",
   "00001001" );    

signal data_aux : std_logic_vector (7 downto 0);
  
begin

reg : process(clk_i, reset_i)
begin
    if reset_i = '0' then
        data_aux <= (Others => '0');
    elsif rising_edge(clk_i) then
        data_aux <= rom(to_integer(unsigned(addr_i)));
    end if;
end process;

data_o <= data_aux;
end Behavioral;
